`timescale 1ns/1ns
`define INV
interface key_expand;

    logic [ 4*4*8 ] round_key_o;
    logic [2:0] current_state;
    logic [ 4*4*8 ] key_in;
    logic [3:0] round;
    logic inv_en;
    logic [3:0] cnt;
    logic rst_n;
    logic clk;

    modport DRV (
        output current_state, key_in, round, cnt, inv_en, rst_n, clk,
        input round_key_o
    );

endinterface //key_expand

class driver;
    virtual key_expand.DRV ke;
    int i, j;
    task run();
        for (i=1 ; i <= 11 ; i = i + 1) begin
            for (j = 0 ; j < 6; j = j + 1) begin
                ke.round <= #5 i;
                ke.cnt <=  #5 j;
                #10;
            end
            $display("%0h\n", ke.round_key_o);
        end
        $finish();
    endtask

endclass

module TB_key_expand;

    // 實例化一個interface
    key_expand ke();

    // 實例化一個driver
    driver drv;

    key_expansion ke_dut(ke.round_key_o, ke.current_state, ke.key_in, ke.round, ke.cnt, ke.inv_en, ke.rst_n, ke.clk);

    event rst_n_reset;

    initial begin
        // Setting Key
        ke.key_in = 128'h2B7E151628AED2A6ABF7158809CF4F3C;
        // ke.key_in = { 8'hBD, 8'h07, 8'hC1, 8'hAC
        //     , 8'h80, 8'h13, 8'h2E, 8'h90
        //     , 8'h16, 8'h19, 8'hF0, 8'h57
        //     , 8'h21, 8'h0B, 8'hA1, 8'h3C };
    end

    initial begin
        ke.current_state <= 3'd1;
        ke.inv_en <= 0;
        ke.clk <= 0;
        ke.rst_n <= 1;
        #10;
        ke.rst_n <= 0;
        #10
        -> rst_n_reset;
        ke.rst_n <= 1;
    end

    always #5 ke.clk <= ~ke.clk;

    initial begin
        drv = new();
        drv.ke = ke;
        wait (rst_n_reset.triggered); 
        #5;
        drv.run();
    end

    initial begin
        $fsdbDumpfile("Key_expand_inv.fsdb");
        $fsdbDumpvars;
        $fsdbDumpMDA();
    end
    
    
endmodule